`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2020/06/04 20:50:03
// Design Name: 
// Module Name: Mux_32
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module Mux_32(
    input SEL,
    input [31:0] in1,
    input [31:0] in2,
    output [31:0] out
    );
    assign out = (SEL)? in2 : in1;
endmodule
